`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 16.12.2024 16:29:58
// Design Name: 
// Module Name: systolicnew
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module systolicnew#(
    parameter WIDTH=16,
    parameter FRAC_BIT=10
)(
input wire clk, 
    input wire rst_n, 
    input wire en, 
    input wire clr,
            input wire                     in_valid,

    input wire signed [WIDTH-1:0] a0, a1, a2,a3,a4,a5,
    input wire signed [WIDTH-1:0] b00, b01, b02, b03, b04, b05,
                                  b10, b11, b12, b13, b14, b15,
                                  b20, b21, b22, b23, b24, b25,
                                  b30, b31, b32, b33, b34, b35,
                                  b40, b41, b42, b43, b44, b45,
                                  b50, b51, b52, b53, b54, b55,   
    output wire signed [WIDTH-1:0] y0, y1,y2,y3,y4,y5,
    output wire                    out_valid,

 wire signed [WIDTH-1:0] y00_in, y01_in, y02_in, y03_in, y04_in, y05_in,

           // *** Valid registers ***
    wire in_valid_reg0, in_valid_reg1, in_valid_reg2, in_valid_reg3, in_valid_reg4, in_valid_reg5, in_valid_reg6, in_valid_reg7, in_valid_reg8, in_valid_reg9, in_valid_reg10, in_valid_reg11, in_valid_reg12,
       a05_out,a15_out,a25_out,a35_out, a45_out, a55_out, // Outputs of systolic array
wire signed [WIDTH-1:0]                                                                                                                                        reg_add_y0out,        
wire signed [WIDTH-1:0]                                                                                                                                        reg50y_1out,                        reg_add_y1out,                        
wire signed [WIDTH-1:0]                                                                                                                                        reg50y_2out,                        reg51y_1out,                        reg_add_y2out,
wire signed [WIDTH-1:0]                                                                                                                                        reg50y_3out,                        reg51y_2out,                        reg52y_1out,                        reg_add_y3out,
wire signed [WIDTH-1:0]                                                                                                                                        reg50y_4out,                        reg51y_3out,                        reg52y_2out,                        reg53y_1out,                        reg_add_y4out,
wire signed [WIDTH-1:0]                                                                                                                                        reg50y_5out,                        reg51y_4out,                        reg52y_3out,                        reg53y_2out,                        reg54y_1out,                         reg_add_y5out,
wire signed [WIDTH-1:0]                                                                                                                                         y50_out,                            y51_out,                            y52_out,                             y53_out,                            y54_out,                            y55_out,
wire signed [WIDTH-1:0]/*reg50*/ reg50_out, /*reg50_1*/ reg50_1out, /*reg50_2*/ reg50_2out, /*reg50_3*/ reg50_3out, /*reg50_4*/ reg50_4out, /*reg50_5*/ a50_in, /*pe50*/ a50_out, /*reg51*/ a51_in, /*pe51*/ a51_out, /*reg52*/ a52_in, /*pe52*/ a52_out, /*reg53*/ a53_in, /*pe53*/ a53_out, /*reg54*/ a54_in, /*pe54*/ a54_out, /*reg55*/ a55_in, /*pe55*/                        
wire signed [WIDTH-1:0]                                                                                                                                        y50_in,                               y51_in,                            y52_in,                             y53_in,                             y54_in,                              y55_in,
wire signed [WIDTH-1:0]                                                                                                                                         y40_out,                            y41_out,                            y42_out,                             y43_out,                            y44_out,                            y45_out,
wire signed [WIDTH-1:0]                        /*reg40*/ reg40_out, /*reg40_1*/ reg40_1out, /*reg40_2*/ reg40_2out, /*reg40_3*/ reg40_3out, /*reg40_4*/ a40_in, /*pe40*/ a40_out, /*reg41*/ a41_in, /*pe41*/ a41_out, /*reg42*/ a42_in, /*pe42*/ a42_out, /*reg43*/ a43_in, /*pe43*/ a43_out, /*reg44*/ a44_in, /*pe44*/ a44_out, /*reg45*/ a45_in, /*pe45*/ 
wire signed [WIDTH-1:0]                                                                                                                                        y40_in,                               y41_in,                            y42_in,                             y43_in,                             y44_in,                              y45_in,
wire signed [WIDTH-1:0]                                                                                                                                         y30_out,                            y31_out,                            y32_out,                             y33_out,                            y34_out,                            y35_out,
wire signed [WIDTH-1:0]                                                /*reg30*/ reg30_out, /*reg30_1*/ reg30_1out, /*reg30_2*/ reg30_2out, /*reg30_3*/ a30_in, /*pe30*/ a30_out, /*reg31*/ a31_in, /*pe31*/ a31_out, /*reg32*/ a32_in, /*pe32*/ a32_out, /*reg33*/ a33_in, /*pe33*/ a33_out, /*reg34*/ a34_in, /*pe34*/ a34_out, /*reg35*/ a35_in, /*pe35*/ 
wire signed [WIDTH-1:0]                                                                                                                                        y30_in,                               y31_in,                            y32_in,                             y33_in,                             y34_in,                              y35_in,
wire signed [WIDTH-1:0]                                                                                                                                         y20_out,                            y21_out,                            y22_out,                             y23_out,                            y24_out,                            y25_out,
wire signed [WIDTH-1:0]                                                                        /*reg20*/ reg20_out, /*reg20_1*/ reg20_1out, /*reg20_2*/ a20_in, /*pe20*/ a20_out, /*reg21*/ a21_in, /*pe21*/ a21_out, /*reg22*/ a22_in, /*pe22*/ a22_out, /*reg23*/ a23_in, /*pe23*/ a23_out, /*reg24*/ a24_in, /*pe24*/ a24_out, /*reg25*/ a25_in, /*pe25*/ 
wire signed [WIDTH-1:0]                                                                                                                                        y20_in,                               y21_in,                            y22_in,                             y23_in,                             y24_in,                              y25_in,
wire signed [WIDTH-1:0]                                                                                                                                         y10_out,                            y11_out,                            y12_out,                             y13_out,                            y14_out,                            y15_out,
wire signed [WIDTH-1:0]                                                                                                /*reg10*/ reg10_out, /*reg10_1*/ a10_in, /*pe10*/ a10_out, /*reg11*/ a11_in, /*pe11*/ a11_out, /*reg12*/ a12_in, /*pe12*/ a12_out, /*reg13*/ a13_in, /*pe13*/ a13_out, /*reg14*/ a14_in, /*pe14*/ a14_out, /*reg15*/ a15_in, /*pe15*/ 
wire signed [WIDTH-1:0]                                                                                                                                        y10_in,                               y11_in,                            y12_in,                             y13_in,                             y14_in,                              y15_in,
wire signed [WIDTH-1:0]                                                                                                                                        y00_out,                            y01_out,                             y02_out,                              y03_out,                            y04_out,                          y05_out,
wire signed [WIDTH-1:0]                                                                                                                       /*reg00*/ a00_in, /*pe00*/ a00_out, /*reg01*/ a01_in, /*pe01*/ a01_out, /*reg02*/ a02_in, /*pe02*/ a02_out, /*reg03*/ a03_in, /*pe03*/ a03_out, /*reg04*/ a04_in, /*pe04*/ a04_out, /*reg05*/ a05_in /*pe05*/ );

    assign y00_in = 0;
    assign y01_in = 0;
    assign y02_in = 0;
    assign y03_in = 0;
    assign y04_in = 0;
    assign y05_in = 0;
    pe #(.WIDTH(WIDTH), .FRAC_BIT(FRAC_BIT)) pe00 (
    .a_in(a00_in),
    .b(b00),
    .y_in(y00_in),
    .a_out(a00_out),
    .y_out(y00_out)
);

pe #(.WIDTH(WIDTH), .FRAC_BIT(FRAC_BIT)) pe01 (
    .a_in(a01_in),
    .b(b01),
    .y_in(y01_in),
    .a_out(a01_out),
    .y_out(y01_out)
);

pe #(.WIDTH(WIDTH), .FRAC_BIT(FRAC_BIT)) pe02 (
    .a_in(a02_in),
    .b(b02),
    .y_in(y02_in),
    .a_out(a02_out),
    .y_out(y02_out)
);

pe #(.WIDTH(WIDTH), .FRAC_BIT(FRAC_BIT)) pe03 (
    .a_in(a03_in),
    .b(b03),
    .y_in(y03_in),
    .a_out(a03_out),
    .y_out(y03_out)
);

pe #(.WIDTH(WIDTH), .FRAC_BIT(FRAC_BIT)) pe04 (
    .a_in(a04_in),
    .b(b04),
    .y_in(y04_in),
    .a_out(a04_out),
    .y_out(y04_out)
);

pe #(.WIDTH(WIDTH), .FRAC_BIT(FRAC_BIT)) pe05 (
    .a_in(a05_in),
    .b(b05),
    .y_in(y05_in),
    .a_out(a05_out),
    .y_out(y05_out)
);

pe #(.WIDTH(WIDTH), .FRAC_BIT(FRAC_BIT)) pe10 (
    .a_in(a10_in),
    .b(b10),
    .y_in(y10_in),
    .a_out(a10_out),
    .y_out(y10_out)
);

pe #(.WIDTH(WIDTH), .FRAC_BIT(FRAC_BIT)) pe11 (
    .a_in(a11_in),
    .b(b11),
    .y_in(y11_in),
    .a_out(a11_out),
    .y_out(y11_out)
);

pe #(.WIDTH(WIDTH), .FRAC_BIT(FRAC_BIT)) pe12 (
    .a_in(a12_in),
    .b(b12),
    .y_in(y12_in),
    .a_out(a12_out),
    .y_out(y12_out)
);

pe #(.WIDTH(WIDTH), .FRAC_BIT(FRAC_BIT)) pe13 (
    .a_in(a13_in),
    .b(b13),
    .y_in(y13_in),
    .a_out(a13_out),
    .y_out(y13_out)
);

pe #(.WIDTH(WIDTH), .FRAC_BIT(FRAC_BIT)) pe14 (
    .a_in(a14_in),
    .b(b14),
    .y_in(y14_in),
    .a_out(a14_out),
    .y_out(y14_out)
);

pe #(.WIDTH(WIDTH), .FRAC_BIT(FRAC_BIT)) pe15 (
    .a_in(a15_in),
    .b(b15),
    .y_in(y15_in),
    .a_out(a15_out),
    .y_out(y15_out)
);

pe #(.WIDTH(WIDTH), .FRAC_BIT(FRAC_BIT)) pe20 (
    .a_in(a20_in),
    .b(b20),
    .y_in(y20_in),
    .a_out(a20_out),
    .y_out(y20_out)
);

pe #(.WIDTH(WIDTH), .FRAC_BIT(FRAC_BIT)) pe21 (
    .a_in(a21_in),
    .b(b21),
    .y_in(y21_in),
    .a_out(a21_out),
    .y_out(y21_out)
);

pe #(.WIDTH(WIDTH), .FRAC_BIT(FRAC_BIT)) pe22 (
    .a_in(a22_in),
    .b(b22),
    .y_in(y22_in),
    .a_out(a22_out),
    .y_out(y22_out)
);

pe #(.WIDTH(WIDTH), .FRAC_BIT(FRAC_BIT)) pe23 (
    .a_in(a23_in),
    .b(b23),
    .y_in(y23_in),
    .a_out(a23_out),
    .y_out(y23_out)
);

pe #(.WIDTH(WIDTH), .FRAC_BIT(FRAC_BIT)) pe24 (
    .a_in(a24_in),
    .b(b24),
    .y_in(y24_in),
    .a_out(a24_out),
    .y_out(y24_out)
);

pe #(.WIDTH(WIDTH), .FRAC_BIT(FRAC_BIT)) pe25 (
    .a_in(a25_in),
    .b(b25),
    .y_in(y25_in),
    .a_out(a25_out),
    .y_out(y25_out)
);

pe #(.WIDTH(WIDTH), .FRAC_BIT(FRAC_BIT)) pe30 (
    .a_in(a30_in),
    .b(b30),
    .y_in(y30_in),
    .a_out(a30_out),
    .y_out(y30_out)
);

pe #(.WIDTH(WIDTH), .FRAC_BIT(FRAC_BIT)) pe31 (
    .a_in(a31_in),
    .b(b31),
    .y_in(y31_in),
    .a_out(a31_out),
    .y_out(y31_out)
);

pe #(.WIDTH(WIDTH), .FRAC_BIT(FRAC_BIT)) pe32 (
    .a_in(a32_in),
    .b(b32),
    .y_in(y32_in),
    .a_out(a32_out),
    .y_out(y32_out)
);

pe #(.WIDTH(WIDTH), .FRAC_BIT(FRAC_BIT)) pe33 (
    .a_in(a33_in),
    .b(b33),
    .y_in(y33_in),
    .a_out(a33_out),
    .y_out(y33_out)
);

pe #(.WIDTH(WIDTH), .FRAC_BIT(FRAC_BIT)) pe34 (
    .a_in(a34_in),
    .b(b34),
    .y_in(y34_in),
    .a_out(a34_out),
    .y_out(y34_out)
);

pe #(.WIDTH(WIDTH), .FRAC_BIT(FRAC_BIT)) pe35 (
    .a_in(a35_in),
    .b(b35),
    .y_in(y35_in),
    .a_out(a35_out),
    .y_out(y35_out)
);

pe #(.WIDTH(WIDTH), .FRAC_BIT(FRAC_BIT)) pe40 (
    .a_in(a40_in),
    .b(b40),
    .y_in(y40_in),
    .a_out(a40_out),
    .y_out(y40_out)
);

pe #(.WIDTH(WIDTH), .FRAC_BIT(FRAC_BIT)) pe41 (
    .a_in(a41_in),
    .b(b41),
    .y_in(y41_in),
    .a_out(a41_out),
    .y_out(y41_out)
);

pe #(.WIDTH(WIDTH), .FRAC_BIT(FRAC_BIT)) pe42 (
    .a_in(a42_in),
    .b(b42),
    .y_in(y42_in),
    .a_out(a42_out),
    .y_out(y42_out)
);

pe #(.WIDTH(WIDTH), .FRAC_BIT(FRAC_BIT)) pe43 (
    .a_in(a43_in),
    .b(b43),
    .y_in(y43_in),
    .a_out(a43_out),
    .y_out(y43_out)
);

pe #(.WIDTH(WIDTH), .FRAC_BIT(FRAC_BIT)) pe44 (
    .a_in(a44_in),
    .b(b44),
    .y_in(y44_in),
    .a_out(a44_out),
    .y_out(y44_out)
);

pe #(.WIDTH(WIDTH), .FRAC_BIT(FRAC_BIT)) pe45 (
    .a_in(a45_in),
    .b(b45),
    .y_in(y45_in),
    .a_out(a45_out),
    .y_out(y45_out)
);

pe #(.WIDTH(WIDTH), .FRAC_BIT(FRAC_BIT)) pe50 (
    .a_in(a50_in),
    .b(b50),
    .y_in(y50_in),
    .a_out(a50_out),
    .y_out(y50_out)
);

pe #(.WIDTH(WIDTH), .FRAC_BIT(FRAC_BIT)) pe51 (
    .a_in(a51_in),
    .b(b51),
    .y_in(y51_in),
    .a_out(a51_out),
    .y_out(y51_out)
);

pe #(.WIDTH(WIDTH), .FRAC_BIT(FRAC_BIT)) pe52 (
    .a_in(a52_in),
    .b(b52),
    .y_in(y52_in),
    .a_out(a52_out),
    .y_out(y52_out)
);

pe #(.WIDTH(WIDTH), .FRAC_BIT(FRAC_BIT)) pe53 (
    .a_in(a53_in),
    .b(b53),
    .y_in(y53_in),
    .a_out(a53_out),
    .y_out(y53_out)
);

pe #(.WIDTH(WIDTH), .FRAC_BIT(FRAC_BIT)) pe54 (
    .a_in(a54_in),
    .b(b54),
    .y_in(y54_in),
    .a_out(a54_out),
    .y_out(y54_out)
);


    pe #(.WIDTH(WIDTH), .FRAC_BIT(FRAC_BIT)) pe55 (
        .a_in(a55_in),
        .b(b55),
        .y_in(y55_in),
        .a_out(a55_out),
        .y_out(y55_out)
    );

    

register #(.WIDTH(WIDTH)) reg00 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(a0),
    .q(a00_in)
);
register #(.WIDTH(WIDTH)) reg01 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(a00_out),
    .q(a01_in)
);
register #(.WIDTH(WIDTH)) reg02 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(a01_out),
    .q(a02_in)
);
register #(.WIDTH(WIDTH)) reg03 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(a02_out),
    .q(a03_in)
);
register #(.WIDTH(WIDTH)) reg04 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(a03_out),
    .q(a04_in)
);
register #(.WIDTH(WIDTH)) reg05 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(a04_out),
    .q(a05_in)
);
register #(.WIDTH(WIDTH)) reg10 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(a1),
    .q(reg10_out)
);

register #(.WIDTH(WIDTH)) reg10_1 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(reg10_out),
    .q(a10_in)
);
register #(.WIDTH(WIDTH)) reg11 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(a10_out),
    .q(a11_in)
);
register #(.WIDTH(WIDTH)) reg12 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(a11_out),
    .q(a12_in)
);
register #(.WIDTH(WIDTH)) reg13 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(a12_out),
    .q(a13_in)
);
register #(.WIDTH(WIDTH)) reg14 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(a13_out),
    .q(a14_in)
);
register #(.WIDTH(WIDTH)) reg15 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(a14_out),
    .q(a15_in)
);
register #(.WIDTH(WIDTH)) reg20 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(a2),
    .q(reg20_out)
);
register #(.WIDTH(WIDTH)) reg20_1 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(reg20_out),
    .q(reg20_1out)
);
register #(.WIDTH(WIDTH)) reg20_2 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(reg20_1out),
    .q(a20_in)
);
register #(.WIDTH(WIDTH)) reg21 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(a20_out),
    .q(a21_in)
);
register #(.WIDTH(WIDTH)) reg22 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(a21_out),
    .q(a22_in)
);
register #(.WIDTH(WIDTH)) reg23 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(a22_out),
    .q(a23_in)
);
register #(.WIDTH(WIDTH)) reg24 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(a23_out),
    .q(a24_in)
);
register #(.WIDTH(WIDTH)) reg25 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(a24_out),
    .q(a25_in)
);
register #(.WIDTH(WIDTH)) reg30 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(a3),
    .q(reg30_out)
);
register #(.WIDTH(WIDTH)) reg30_1 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(reg30_out),
    .q(reg30_1out)
);
register #(.WIDTH(WIDTH)) reg30_2 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(reg30_1out),
    .q(reg30_2out)
);
register #(.WIDTH(WIDTH)) reg30_3 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(reg30_2out),
    .q(a30_in)
);
register #(.WIDTH(WIDTH)) reg31 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(a30_out),
    .q(a31_in)
);
register #(.WIDTH(WIDTH)) reg32 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(a31_out),
    .q(a32_in)
);
register #(.WIDTH(WIDTH)) reg33 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(a32_out),
    .q(a33_in)
);
register #(.WIDTH(WIDTH)) reg34 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(a33_out),
    .q(a34_in)
);
register #(.WIDTH(WIDTH)) reg35 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(a34_out),
    .q(a35_in)
);
register #(.WIDTH(WIDTH)) reg40 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(a4),
    .q(reg40_out)
);
register #(.WIDTH(WIDTH)) reg40_1 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(reg40_out),
    .q(reg40_1out)
);
register #(.WIDTH(WIDTH)) reg40_2 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(reg40_1out),
    .q(reg40_2out)
);
register #(.WIDTH(WIDTH)) reg40_3 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(reg40_2out),
    .q(reg40_3out)
);
register #(.WIDTH(WIDTH)) reg40_4 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(reg40_3out),
    .q(a40_in)
);

register #(.WIDTH(WIDTH)) reg41 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(a40_out),
    .q(a41_in)
);
register #(.WIDTH(WIDTH)) reg42 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(a41_out),
    .q(a42_in)
);
register #(.WIDTH(WIDTH)) reg43 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(a42_out),
    .q(a43_in)
);
register #(.WIDTH(WIDTH)) reg44 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(a43_out),
    .q(a44_in)
);
register #(.WIDTH(WIDTH)) reg45 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(a44_out),
    .q(a45_in)
);
register #(.WIDTH(WIDTH)) reg50 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(a5),
    .q(reg50_out)
);
register #(.WIDTH(WIDTH)) reg50_1 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(reg50_out),
    .q(reg50_1out)
);
register #(.WIDTH(WIDTH)) reg50_2 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(reg50_1out),
    .q(reg50_2out)
);
register #(.WIDTH(WIDTH)) reg50_3 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(reg50_2out),
    .q(reg50_3out)
);
register #(.WIDTH(WIDTH)) reg50_4 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(reg50_3out),
    .q(reg50_4out)
);
register #(.WIDTH(WIDTH)) reg50_5 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(reg50_4out),
    .q(a50_in)
);
register #(.WIDTH(WIDTH)) reg51 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(a50_out),
    .q(a51_in)
);
register #(.WIDTH(WIDTH)) reg52 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(a51_out),
    .q(a52_in)
);
register #(.WIDTH(WIDTH)) reg53 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(a52_out),
    .q(a53_in)
);
register #(.WIDTH(WIDTH)) reg54 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(a53_out),
    .q(a54_in)
);
register #(.WIDTH(WIDTH)) reg55 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(a54_out),
    .q(a55_in)
);

register #(.WIDTH(WIDTH)) reg00y (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(y00_out),
    .q(y10_in)
);
register #(.WIDTH(WIDTH)) reg01y (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(y01_out),
    .q(y11_in)
);
register #(.WIDTH(WIDTH)) reg02y (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(y02_out),
    .q(y12_in)
);
register #(.WIDTH(WIDTH)) reg03y (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(y03_out),
    .q(y13_in)
);
register #(.WIDTH(WIDTH)) reg04y (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(y04_out),
    .q(y14_in)
);
register #(.WIDTH(WIDTH)) reg05y (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(y05_out),
    .q(y15_in)
);
register #(.WIDTH(WIDTH)) reg10y (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(y10_out),
    .q(y20_in)
);
register #(.WIDTH(WIDTH)) reg11y (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(y11_out),
    .q(y21_in)
);
register #(.WIDTH(WIDTH)) reg12y (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(y12_out),
    .q(y22_in)
);
register #(.WIDTH(WIDTH)) reg13y (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(y13_out),
    .q(y23_in)
);
register #(.WIDTH(WIDTH)) reg14y (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(y14_out),
    .q(y24_in)
);
register #(.WIDTH(WIDTH)) reg15y (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(y15_out),
    .q(y25_in)
);
register #(.WIDTH(WIDTH)) reg20y (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(y20_out),
    .q(y30_in)
);
register #(.WIDTH(WIDTH)) reg21y (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(y21_out),
    .q(y31_in)
);
register #(.WIDTH(WIDTH)) reg22y (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(y22_out),
    .q(y32_in)
);
register #(.WIDTH(WIDTH)) reg23y (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(y23_out),
    .q(y33_in)
);
register #(.WIDTH(WIDTH)) reg24y (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(y24_out),
    .q(y34_in)
);
register #(.WIDTH(WIDTH)) reg25y (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(y25_out),
    .q(y35_in)
);
register #(.WIDTH(WIDTH)) reg30y (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(y30_out),
    .q(y40_in)
);
register #(.WIDTH(WIDTH)) reg31y (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(y31_out),
    .q(y41_in)
);
register #(.WIDTH(WIDTH)) reg32y (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(y32_out),
    .q(y42_in)
);
register #(.WIDTH(WIDTH)) reg33y (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(y33_out),
    .q(y43_in)
);
register #(.WIDTH(WIDTH)) reg34y (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(y34_out),
    .q(y44_in)
);
register #(.WIDTH(WIDTH)) reg35y (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(y35_out),
    .q(y45_in)
);
register #(.WIDTH(WIDTH)) reg40y (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(y40_out),
    .q(y50_in)
);
register #(.WIDTH(WIDTH)) reg41y (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(y41_out),
    .q(y51_in)
);
register #(.WIDTH(WIDTH)) reg42y (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(y42_out),
    .q(y52_in)
);
register #(.WIDTH(WIDTH)) reg43y (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(y43_out),
    .q(y53_in)
);
register #(.WIDTH(WIDTH)) reg44y (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(y44_out),
    .q(y54_in)
);
register #(.WIDTH(WIDTH)) reg45y (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(y45_out),
    .q(y55_in)
);
register #(.WIDTH(WIDTH)) reg50y (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(reg50y_1out),
    .q(reg_add_y0out)
);
register #(.WIDTH(WIDTH)) reg50y_1 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(reg50y_2out),
    .q(reg50y_1out)
);
register #(.WIDTH(WIDTH)) reg50y_2 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(reg50y_3out),
    .q(reg50y_2out)
);
register #(.WIDTH(WIDTH)) reg50y_3 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(reg50y_4out),
    .q(reg50y_3out)
);
register #(.WIDTH(WIDTH)) reg50y_4 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(reg50y_5out),
    .q(reg50y_4out)
);
register #(.WIDTH(WIDTH)) reg50y_5 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(y50_out),
    .q(reg50y_5out)
);
register #(.WIDTH(WIDTH)) reg51y (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(reg51y_1out),
    .q(reg_add_y1out)
);
register #(.WIDTH(WIDTH)) reg51y_1 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(reg51y_2out),
    .q(reg51y_1out)
);
register #(.WIDTH(WIDTH)) reg51y_2 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(reg51y_3out),
    .q(reg51y_2out)
);
register #(.WIDTH(WIDTH)) reg51y_3 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(reg51y_4out),
    .q(reg51y_3out)
);
register #(.WIDTH(WIDTH)) reg51y_4 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(y51_out),
    .q(reg51y_4out)
);
register #(.WIDTH(WIDTH)) reg52y (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(reg52y_1out),
    .q(reg_add_y2out)
);
register #(.WIDTH(WIDTH)) reg52y_1 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(reg52y_2out),
    .q(reg52y_1out)
);
register #(.WIDTH(WIDTH)) reg52y_2 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(reg52y_3out),
    .q(reg52y_2out)
);
register #(.WIDTH(WIDTH)) reg52y_3 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(y52_out),
    .q(reg52y_3out)
);

register #(.WIDTH(WIDTH)) reg53y (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(reg53y_1out),
    .q(reg_add_y3out)
);
register #(.WIDTH(WIDTH)) reg53y_1 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(reg53y_2out),
    .q(reg53y_1out)
);
register #(.WIDTH(WIDTH)) reg53y_2 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(y53_out),
    .q(reg53y_2out)
);

register #(.WIDTH(WIDTH)) reg54y (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(reg54y_1out),
    .q(reg_add_y4out)
);
register #(.WIDTH(WIDTH)) reg54y_1 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(y54_out),
    .q(reg54y_1out)
);

register #(.WIDTH(WIDTH)) reg55y (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(y55_out),
    .q(reg_add_y5out)
);

// ADDITIONAL TIMING ADJUST REGISTER FOR OUTPUT
register #(.WIDTH(WIDTH)) reg_add_y0 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(reg_add_y0out),
    .q(y0)
);
register #(.WIDTH(WIDTH)) reg_add_y1 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(reg_add_y1out),
    .q(y1)
);
register #(.WIDTH(WIDTH)) reg_add_y2 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(reg_add_y2out),
    .q(y2)
);
register #(.WIDTH(WIDTH)) reg_add_y3 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(reg_add_y3out),
    .q(y3)
);
register #(.WIDTH(WIDTH)) reg_add_y4 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(reg_add_y4out),
    .q(y4)
);
register #(.WIDTH(WIDTH)) reg_add_y5 (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .clr(clr),
    .d(reg_add_y0out),
    .q(y5)
);
   // *** Valid registers ***
    register #(1) reg_valid_0(clk, rst_n, en, clr, in_valid,      in_valid_reg0); 
    register #(1) reg_valid_1(clk, rst_n, en, clr, in_valid_reg0, in_valid_reg1);
    register #(1) reg_valid_2(clk, rst_n, en, clr, in_valid_reg1, in_valid_reg2);
    register #(1) reg_valid_3(clk, rst_n, en, clr, in_valid_reg2, in_valid_reg3);
    register #(1) reg_valid_4(clk, rst_n, en, clr, in_valid_reg3, in_valid_reg4);
    register #(1) reg_valid_5(clk, rst_n, en, clr, in_valid_reg4, in_valid_reg5);
    register #(1) reg_valid_6(clk, rst_n, en, clr, in_valid_reg5, in_valid_reg6);
    register #(1) reg_valid_7(clk, rst_n, en, clr, in_valid_reg6, in_valid_reg7);
    register #(1) reg_valid_8(clk, rst_n, en, clr, in_valid_reg7, in_valid_reg8);
    register #(1) reg_valid_9(clk, rst_n, en, clr, in_valid_reg8, in_valid_reg9);
    register #(1) reg_valid_10(clk, rst_n, en, clr, in_valid_reg9, in_valid_reg10);
    register #(1) reg_valid_11(clk, rst_n, en, clr, in_valid_reg10, in_valid_reg11);    
    register #(1) reg_valid_12(clk, rst_n, en, clr, in_valid_reg11, in_valid_reg12);  
    assign out_valid = in_valid_reg12;


endmodule
